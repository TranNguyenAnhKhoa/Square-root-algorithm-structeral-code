`timescale 1ps/1ps
module tb_sra();


endmodule

